library verilog;
use verilog.vl_types.all;
entity top is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        A1              : in     vl_logic;
        SW_choose       : in     vl_logic;
        SW1             : in     vl_logic;
        SW2             : in     vl_logic;
        D               : in     vl_logic_vector(7 downto 0);
        addr            : out    vl_logic_vector(15 downto 0);
        rambus          : out    vl_logic_vector(7 downto 0);
        data            : out    vl_logic_vector(7 downto 0);
        HEX0            : out    vl_logic_vector(6 downto 0);
        HEX1            : out    vl_logic_vector(6 downto 0);
        HEX2            : out    vl_logic_vector(6 downto 0);
        HEX3            : out    vl_logic_vector(6 downto 0);
        HEX4            : out    vl_logic_vector(6 downto 0);
        HEX5            : out    vl_logic_vector(6 downto 0);
        HEX6            : out    vl_logic_vector(6 downto 0);
        HEX7            : out    vl_logic_vector(6 downto 0);
        acdbus          : out    vl_logic_vector(7 downto 0);
        rdbus           : out    vl_logic_vector(7 downto 0);
        cpustate_led    : out    vl_logic_vector(1 downto 0);
        check_out       : out    vl_logic_vector(7 downto 0);
        quick_low_led   : out    vl_logic;
        read_led        : out    vl_logic;
        write_led       : out    vl_logic;
        arload_led      : out    vl_logic;
        pcinc_led       : out    vl_logic;
        pcload_led      : out    vl_logic;
        drload_led      : out    vl_logic;
        trload_led      : out    vl_logic;
        irload_led      : out    vl_logic;
        rload_led       : out    vl_logic;
        acload_led      : out    vl_logic;
        zload_led       : out    vl_logic;
        pcbus_led       : out    vl_logic;
        drhbus_led      : out    vl_logic;
        drlbus_led      : out    vl_logic;
        trbus_led       : out    vl_logic;
        rbus_led        : out    vl_logic;
        acbus_led       : out    vl_logic;
        membus_led      : out    vl_logic;
        irbus_led       : out    vl_logic;
        busmem_led      : out    vl_logic;
        clr_led         : out    vl_logic
    );
end top;
